/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module CC_SCREENCOMPARATOR (
//////////// OUTPUTS //////////
	CC_SCREENCOMPARATOR_0,
	CC_SCREENCOMPARATOR_1,
	CC_SCREENCOMPARATOR_2,
	CC_SCREENCOMPARATOR_3,
	CC_SCREENCOMPARATOR_4,
	CC_SCREENCOMPARATOR_5,
	CC_SCREENCOMPARATOR_6,
	CC_SCREENCOMPARATOR_7,
//////////// INPUTS //////////
	CC_SCREENCOMPARATOR_POINT_0,
	CC_SCREENCOMPARATOR_POINT_1,
	CC_SCREENCOMPARATOR_POINT_2,
	CC_SCREENCOMPARATOR_POINT_3,
	CC_SCREENCOMPARATOR_POINT_4,
	CC_SCREENCOMPARATOR_POINT_5,
	CC_SCREENCOMPARATOR_POINT_6,
	CC_SCREENCOMPARATOR_POINT_7,
	CC_SCREENCOMPARATOR_POINT_8,
	CC_SCREENCOMPARATOR_POINT_9,
	CC_SCREENCOMPARATOR_POINT_10,
	CC_SCREENCOMPARATOR_POINT_11,
	CC_SCREENCOMPARATOR_POINT_12,
	CC_SCREENCOMPARATOR_POINT_13,
	CC_SCREENCOMPARATOR_POINT_14,
	
	CC_SCREENCOMPARATOR_BACK_0,
	CC_SCREENCOMPARATOR_BACK_1,
	CC_SCREENCOMPARATOR_BACK_2,
	CC_SCREENCOMPARATOR_BACK_3,
	CC_SCREENCOMPARATOR_BACK_4,
	CC_SCREENCOMPARATOR_BACK_5,
	CC_SCREENCOMPARATOR_BACK_6,
	CC_SCREENCOMPARATOR_BACK_7,
	CC_SCREENCOMPARATOR_BACK_8,
	CC_SCREENCOMPARATOR_BACK_9,
	CC_SCREENCOMPARATOR_BACK_10,
	CC_SCREENCOMPARATOR_BACK_11,
	CC_SCREENCOMPARATOR_BACK_12,
	CC_SCREENCOMPARATOR_BACK_13,
	CC_SCREENCOMPARATOR_BACK_14,
	
	CC_SCREENCOMPARATOR_LOSE_0,
	CC_SCREENCOMPARATOR_LOSE_1,
	CC_SCREENCOMPARATOR_LOSE_2,
	CC_SCREENCOMPARATOR_LOSE_3,
	CC_SCREENCOMPARATOR_LOSE_4,
	CC_SCREENCOMPARATOR_LOSE_5,
	CC_SCREENCOMPARATOR_LOSE_6,
	CC_SCREENCOMPARATOR_LOSE_7,
	
	CC_SCREENCOMPARATOR_WIN_0,
	CC_SCREENCOMPARATOR_WIN_1,
	CC_SCREENCOMPARATOR_WIN_2,
	CC_SCREENCOMPARATOR_WIN_3,
	CC_SCREENCOMPARATOR_WIN_4,
	CC_SCREENCOMPARATOR_WIN_5,
	CC_SCREENCOMPARATOR_WIN_6,
	CC_SCREENCOMPARATOR_WIN_7,
	
	CC_SCREENCOMPARATOR_LOSE,
	CC_SCREENCOMPARATOR_WIN
);
//=======================================================
//  PORT declarations
//=======================================================
output reg [7:0]CC_SCREENCOMPARATOR_0;
output reg [7:0]CC_SCREENCOMPARATOR_1;
output reg [7:0]CC_SCREENCOMPARATOR_2;
output reg [7:0]CC_SCREENCOMPARATOR_3;
output reg [7:0]CC_SCREENCOMPARATOR_4;
output reg [7:0]CC_SCREENCOMPARATOR_5;
output reg [7:0]CC_SCREENCOMPARATOR_6;
output reg [7:0]CC_SCREENCOMPARATOR_7;

input [7:0]CC_SCREENCOMPARATOR_POINT_0;
input [7:0]CC_SCREENCOMPARATOR_POINT_1;
input [7:0]CC_SCREENCOMPARATOR_POINT_2;
input [7:0]CC_SCREENCOMPARATOR_POINT_3;
input [7:0]CC_SCREENCOMPARATOR_POINT_4;
input [7:0]CC_SCREENCOMPARATOR_POINT_5;
input [7:0]CC_SCREENCOMPARATOR_POINT_6;
input [7:0]CC_SCREENCOMPARATOR_POINT_7;
input [7:0]CC_SCREENCOMPARATOR_POINT_8;
input [7:0]CC_SCREENCOMPARATOR_POINT_9;
input [7:0]CC_SCREENCOMPARATOR_POINT_10;
input [7:0]CC_SCREENCOMPARATOR_POINT_11;
input [7:0]CC_SCREENCOMPARATOR_POINT_12;
input [7:0]CC_SCREENCOMPARATOR_POINT_13;
input [7:0]CC_SCREENCOMPARATOR_POINT_14;

input	[7:0]CC_SCREENCOMPARATOR_BACK_0;
input	[7:0]CC_SCREENCOMPARATOR_BACK_1;
input	[7:0]CC_SCREENCOMPARATOR_BACK_2;
input	[7:0]CC_SCREENCOMPARATOR_BACK_3;
input	[7:0]CC_SCREENCOMPARATOR_BACK_4;
input	[7:0]CC_SCREENCOMPARATOR_BACK_5;
input	[7:0]CC_SCREENCOMPARATOR_BACK_6;
input	[7:0]CC_SCREENCOMPARATOR_BACK_7;
input	[7:0]CC_SCREENCOMPARATOR_BACK_8;
input	[7:0]CC_SCREENCOMPARATOR_BACK_9;
input	[7:0]CC_SCREENCOMPARATOR_BACK_10;
input	[7:0]CC_SCREENCOMPARATOR_BACK_11;
input	[7:0]CC_SCREENCOMPARATOR_BACK_12;
input	[7:0]CC_SCREENCOMPARATOR_BACK_13;
input	[7:0]CC_SCREENCOMPARATOR_BACK_14;
	
input [7:0]CC_SCREENCOMPARATOR_LOSE_0;
input [7:0]CC_SCREENCOMPARATOR_LOSE_1;
input [7:0]CC_SCREENCOMPARATOR_LOSE_2;
input [7:0]CC_SCREENCOMPARATOR_LOSE_3;
input [7:0]CC_SCREENCOMPARATOR_LOSE_4;
input [7:0]CC_SCREENCOMPARATOR_LOSE_5;
input [7:0]CC_SCREENCOMPARATOR_LOSE_6;
input [7:0]CC_SCREENCOMPARATOR_LOSE_7;

input [7:0]CC_SCREENCOMPARATOR_WIN_0;
input [7:0]CC_SCREENCOMPARATOR_WIN_1;
input [7:0]CC_SCREENCOMPARATOR_WIN_2;
input [7:0]CC_SCREENCOMPARATOR_WIN_3;
input [7:0]CC_SCREENCOMPARATOR_WIN_4;
input [7:0]CC_SCREENCOMPARATOR_WIN_5;
input [7:0]CC_SCREENCOMPARATOR_WIN_6;
input [7:0]CC_SCREENCOMPARATOR_WIN_7;

input [2:0]CC_SCREENCOMPARATOR_LOSE;
input	[3:0]CC_SCREENCOMPARATOR_WIN;
//=======================================================
//  Structural coding
//=======================================================
always @(*)
begin
	if (CC_SCREENCOMPARATOR_LOSE == 2'b10)
		begin
		CC_SCREENCOMPARATOR_0 = CC_SCREENCOMPARATOR_LOSE_0;
		CC_SCREENCOMPARATOR_1 = CC_SCREENCOMPARATOR_LOSE_1;
		CC_SCREENCOMPARATOR_2 = CC_SCREENCOMPARATOR_LOSE_2;
		CC_SCREENCOMPARATOR_3 = CC_SCREENCOMPARATOR_LOSE_3;
		CC_SCREENCOMPARATOR_4 = CC_SCREENCOMPARATOR_LOSE_4;
		CC_SCREENCOMPARATOR_5 = CC_SCREENCOMPARATOR_LOSE_5;
		CC_SCREENCOMPARATOR_6 = CC_SCREENCOMPARATOR_LOSE_6;
		CC_SCREENCOMPARATOR_7 = CC_SCREENCOMPARATOR_LOSE_7;
		end
	else if (CC_SCREENCOMPARATOR_WIN == 2'b11)
		begin
		CC_SCREENCOMPARATOR_0 = CC_SCREENCOMPARATOR_WIN_0;
		CC_SCREENCOMPARATOR_1 = CC_SCREENCOMPARATOR_WIN_1;
		CC_SCREENCOMPARATOR_2 = CC_SCREENCOMPARATOR_WIN_2;
		CC_SCREENCOMPARATOR_3 = CC_SCREENCOMPARATOR_WIN_3;
		CC_SCREENCOMPARATOR_4 = CC_SCREENCOMPARATOR_WIN_4;
		CC_SCREENCOMPARATOR_5 = CC_SCREENCOMPARATOR_WIN_5;
		CC_SCREENCOMPARATOR_6 = CC_SCREENCOMPARATOR_WIN_6;
		CC_SCREENCOMPARATOR_7 = CC_SCREENCOMPARATOR_WIN_7;
		end
	else if ((CC_SCREENCOMPARATOR_POINT_7 | CC_SCREENCOMPARATOR_POINT_8 | CC_SCREENCOMPARATOR_POINT_9 | CC_SCREENCOMPARATOR_POINT_10 | CC_SCREENCOMPARATOR_POINT_11 | CC_SCREENCOMPARATOR_POINT_12 | CC_SCREENCOMPARATOR_POINT_13 | CC_SCREENCOMPARATOR_POINT_14) != 8'b00000000)
		begin
		CC_SCREENCOMPARATOR_0 = CC_SCREENCOMPARATOR_BACK_7 | CC_SCREENCOMPARATOR_POINT_7;
		CC_SCREENCOMPARATOR_1 = CC_SCREENCOMPARATOR_BACK_8 | CC_SCREENCOMPARATOR_POINT_8;
		CC_SCREENCOMPARATOR_2 = CC_SCREENCOMPARATOR_BACK_9 | CC_SCREENCOMPARATOR_POINT_9;
		CC_SCREENCOMPARATOR_3 = CC_SCREENCOMPARATOR_BACK_10 | CC_SCREENCOMPARATOR_POINT_10;
		CC_SCREENCOMPARATOR_4 = CC_SCREENCOMPARATOR_BACK_11 | CC_SCREENCOMPARATOR_POINT_11;
		CC_SCREENCOMPARATOR_5 = CC_SCREENCOMPARATOR_BACK_12 | CC_SCREENCOMPARATOR_POINT_12;
		CC_SCREENCOMPARATOR_6 = CC_SCREENCOMPARATOR_BACK_13 | CC_SCREENCOMPARATOR_POINT_13;
		CC_SCREENCOMPARATOR_7 = CC_SCREENCOMPARATOR_BACK_14 | CC_SCREENCOMPARATOR_POINT_14;
		end
	else
		begin
		CC_SCREENCOMPARATOR_0 = CC_SCREENCOMPARATOR_BACK_0 | CC_SCREENCOMPARATOR_POINT_0;
		CC_SCREENCOMPARATOR_1 = CC_SCREENCOMPARATOR_BACK_1 | CC_SCREENCOMPARATOR_POINT_1;
		CC_SCREENCOMPARATOR_2 = CC_SCREENCOMPARATOR_BACK_2 | CC_SCREENCOMPARATOR_POINT_2;
		CC_SCREENCOMPARATOR_3 = CC_SCREENCOMPARATOR_BACK_3 | CC_SCREENCOMPARATOR_POINT_3;
		CC_SCREENCOMPARATOR_4 = CC_SCREENCOMPARATOR_BACK_4 | CC_SCREENCOMPARATOR_POINT_4;
		CC_SCREENCOMPARATOR_5 = CC_SCREENCOMPARATOR_BACK_5 | CC_SCREENCOMPARATOR_POINT_5;
		CC_SCREENCOMPARATOR_6 = CC_SCREENCOMPARATOR_BACK_6 | CC_SCREENCOMPARATOR_POINT_6;
		CC_SCREENCOMPARATOR_7 = CC_SCREENCOMPARATOR_BACK_7 | CC_SCREENCOMPARATOR_POINT_7;
		end
end

endmodule

