/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module CC_COLLISIONCOMPARATOR (
//////////// OUTPUTS //////////
	CC_COLLISIONCOMPARATOR_EXIT,
//////////// INPUTS //////////
	CC_COLLISIONCOMPARATOR_POINT_0,
	CC_COLLISIONCOMPARATOR_POINT_1,
	CC_COLLISIONCOMPARATOR_POINT_2,
	CC_COLLISIONCOMPARATOR_POINT_3,
	CC_COLLISIONCOMPARATOR_POINT_4,
	CC_COLLISIONCOMPARATOR_POINT_5,
	CC_COLLISIONCOMPARATOR_POINT_6,
	CC_COLLISIONCOMPARATOR_POINT_7,
	CC_COLLISIONCOMPARATOR_POINT_8,
	CC_COLLISIONCOMPARATOR_POINT_9,
	CC_COLLISIONCOMPARATOR_POINT_10,
	CC_COLLISIONCOMPARATOR_POINT_11,
	CC_COLLISIONCOMPARATOR_POINT_12,
	CC_COLLISIONCOMPARATOR_POINT_13,
	CC_COLLISIONCOMPARATOR_POINT_14,
	
	CC_COLLISIONCOMPARATOR_BACK_0,
	CC_COLLISIONCOMPARATOR_BACK_1,
	CC_COLLISIONCOMPARATOR_BACK_2,
	CC_COLLISIONCOMPARATOR_BACK_3,
	CC_COLLISIONCOMPARATOR_BACK_4,
	CC_COLLISIONCOMPARATOR_BACK_5,
	CC_COLLISIONCOMPARATOR_BACK_6,
	CC_COLLISIONCOMPARATOR_BACK_7,
	CC_COLLISIONCOMPARATOR_BACK_8,
	CC_COLLISIONCOMPARATOR_BACK_9,
	CC_COLLISIONCOMPARATOR_BACK_10,
	CC_COLLISIONCOMPARATOR_BACK_11,
	CC_COLLISIONCOMPARATOR_BACK_12,
	CC_COLLISIONCOMPARATOR_BACK_13,
	CC_COLLISIONCOMPARATOR_BACK_14,
	CC_COLLISIONCOMPARATOR_LOSE,
	CC_COLLISIONCOMPARATOR_WIN
);
//=======================================================
//  PORT declarations
//=======================================================
output reg CC_COLLISIONCOMPARATOR_EXIT;

input [7:0]CC_COLLISIONCOMPARATOR_POINT_0;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_1;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_2;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_3;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_4;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_5;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_6;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_7;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_8;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_9;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_10;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_11;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_12;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_13;
input [7:0]CC_COLLISIONCOMPARATOR_POINT_14;
	
input [7:0]CC_COLLISIONCOMPARATOR_BACK_0;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_1;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_2;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_3;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_4;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_5;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_6;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_7;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_8;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_9;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_10;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_11;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_12;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_13;
input [7:0]CC_COLLISIONCOMPARATOR_BACK_14;
input	[2:0]CC_COLLISIONCOMPARATOR_LOSE;
input	[3:0]CC_COLLISIONCOMPARATOR_WIN;
//=======================================================
//  Structural coding
//=======================================================
always @(*)
begin
	if (CC_COLLISIONCOMPARATOR_LOSE == 2'b10)
		CC_COLLISIONCOMPARATOR_EXIT = 1'b0;
	else if (CC_COLLISIONCOMPARATOR_WIN == 2'b11)
		CC_COLLISIONCOMPARATOR_EXIT = 1'b0;
	else if((CC_COLLISIONCOMPARATOR_BACK_0 & CC_COLLISIONCOMPARATOR_POINT_0 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_1 & CC_COLLISIONCOMPARATOR_POINT_1 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_2 & CC_COLLISIONCOMPARATOR_POINT_2 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_3 & CC_COLLISIONCOMPARATOR_POINT_3 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_4 & CC_COLLISIONCOMPARATOR_POINT_4 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_5 & CC_COLLISIONCOMPARATOR_POINT_5 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_6 & CC_COLLISIONCOMPARATOR_POINT_6 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_7 & CC_COLLISIONCOMPARATOR_POINT_7 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_8 & CC_COLLISIONCOMPARATOR_POINT_8 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_9 & CC_COLLISIONCOMPARATOR_POINT_9 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_10 & CC_COLLISIONCOMPARATOR_POINT_10 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_11 & CC_COLLISIONCOMPARATOR_POINT_11 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_12 & CC_COLLISIONCOMPARATOR_POINT_12 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_13 & CC_COLLISIONCOMPARATOR_POINT_13 != 8'b00000000) || (CC_COLLISIONCOMPARATOR_BACK_14 & CC_COLLISIONCOMPARATOR_POINT_14 != 8'b00000000))
		CC_COLLISIONCOMPARATOR_EXIT = 1'b1;
	else 
		CC_COLLISIONCOMPARATOR_EXIT = 1'b0;
end

endmodule

