/*######################################################################
//#	G0B1T: HDL EXAMPLES. 2018.
//######################################################################
//# Copyright (C) 2018. F.E.Segura-Quijano (FES) fsegura@uniandes.edu.co
//# 
//# This program is free software: you can redistribute it and/or modify
//# it under the terms of the GNU General Public License as published by
//# the Free Software Foundation, version 3 of the License.
//#
//# This program is distributed in the hope that it will be useful,
//# but WITHOUT ANY WARRANTY; without even the implied warranty of
//# MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//# GNU General Public License for more details.
//#
//# You should have received a copy of the GNU General Public License
//# along with this program.  If not, see <http://www.gnu.org/licenses/>
//####################################################################*/
//=======================================================
//  MODULE Definition
//=======================================================
module BB_SYSTEM (
//////////// OUTPUTS //////////
	BB_SYSTEM_display_OutBUS,
	BB_SYSTEM_max7219DIN_Out,
	BB_SYSTEM_max7219NCS_Out,
	BB_SYSTEM_max7219CLK_Out,

	BB_SYSTEM_startButton_Out, 
	BB_SYSTEM_upButton_Out,
	BB_SYSTEM_downButton_Out,
	BB_SYSTEM_leftButton_Out,
	BB_SYSTEM_rightButton_Out,
	BB_SYSTEM_TEST0,
	BB_SYSTEM_TEST1,
	BB_SYSTEM_TEST2,

//////////// INPUTS //////////
	BB_SYSTEM_CLOCK_50,
	BB_SYSTEM_RESET_InHigh,
	BB_SYSTEM_startButton_InLow, 
	BB_SYSTEM_upButton_InLow,
	BB_SYSTEM_downButton_InLow,
	BB_SYSTEM_leftButton_InLow,
	BB_SYSTEM_rightButton_InLow
);
//=======================================================
//  PARAMETER declarations
//=======================================================
 parameter DATAWIDTH_BUS = 8;
 parameter PRESCALER_DATAWIDTH = 23;
 parameter DISPLAY_DATAWIDTH = 12;
 
 parameter DATA_FIXED_INITREGPOINT_14 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_13 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_12 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_11 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_10 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_9 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_8 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_7 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_6 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_5 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_4 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_3 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_2 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_1 = 8'b00000000;
 parameter DATA_FIXED_INITREGPOINT_0 = 8'b00010000;
 
 parameter DATA_FIXED_INITREGBACKG_14 = 8'b11100111;
 
 parameter INITREGBACKG_13 = 8'b00000000;
 parameter INITREGBACKG_12 = 8'b00111000;
 parameter INITREGBACKG_11 = 8'b00000000;
 parameter INITREGBACKG_10 = 8'b11001100;
 parameter INITREGBACKG_9 = 8'b00000000;
 parameter INITREGBACKG_8 = 8'b01110000;
 parameter INITREGBACKG_7 = 8'b00000000;
 parameter INITREGBACKG_6 = 8'b00001110;
 parameter INITREGBACKG_5 = 8'b00000000;
 parameter INITREGBACKG_4 = 8'b00111000;
 parameter INITREGBACKG_3 = 8'b00000000;
 parameter INITREGBACKG_2 = 8'b11100000;
 parameter INITREGBACKG_1 = 8'b00000000;
 parameter INITREGBACKG_0 = 8'b00000000;
 
 parameter INITREGBACKG_13_1 = 8'b00000000;
 parameter INITREGBACKG_12_1 = 8'b00011110;
 parameter INITREGBACKG_11_1 = 8'b00000000;
 parameter INITREGBACKG_10_1 = 8'b11100111;
 parameter INITREGBACKG_9_1 = 8'b11100111;
 parameter INITREGBACKG_8_1 = 8'b00000000;
 parameter INITREGBACKG_7_1 = 8'b00000000;
 parameter INITREGBACKG_6_1 = 8'b00111000;
 parameter INITREGBACKG_5_1 = 8'b00000000;
 parameter INITREGBACKG_4_1 = 8'b11101110;
 parameter INITREGBACKG_3_1 = 8'b00000000;
 parameter INITREGBACKG_2_1 = 8'b11110000;
 parameter INITREGBACKG_1_1 = 8'b00000000;
 parameter INITREGBACKG_0_1 = 8'b00000000;
 
 parameter INITREGBACKG_13_2 = 8'b00000000;
 parameter INITREGBACKG_12_2 = 8'b11100000;
 parameter INITREGBACKG_11_2 = 8'b00000000;
 parameter INITREGBACKG_10_2 = 8'b11000110;
 parameter INITREGBACKG_9_2 = 8'b11100000;
 parameter INITREGBACKG_8_2 = 8'b00011100;
 parameter INITREGBACKG_7_2 = 8'b00000000;
 parameter INITREGBACKG_6_2 = 8'b00111000;
 parameter INITREGBACKG_5_2 = 8'b00000000;
 parameter INITREGBACKG_4_2 = 8'b11011111;
 parameter INITREGBACKG_3_2 = 8'b11000111;
 parameter INITREGBACKG_2_2 = 8'b11100111;
 parameter INITREGBACKG_1_2 = 8'b00000000;
 parameter INITREGBACKG_0_2 = 8'b00000000;
 
 parameter INITREGBACKG_13_3 = 8'b00000000;
 parameter INITREGBACKG_12_3 = 8'b01110000;
 parameter INITREGBACKG_11_3 = 8'b00000000;
 parameter INITREGBACKG_10_3 = 8'b10101010;
 parameter INITREGBACKG_9_3 = 8'b01110000;
 parameter INITREGBACKG_8_3 = 8'b00001110;
 parameter INITREGBACKG_7_3 = 8'b00000000;
 parameter INITREGBACKG_6_3 = 8'b00111100;
 parameter INITREGBACKG_5_3 = 8'b00000000;
 parameter INITREGBACKG_4_3 = 8'b11100111;
 parameter INITREGBACKG_3_3 = 8'b11100111;
 parameter INITREGBACKG_2_3 = 8'b11100111;
 parameter INITREGBACKG_1_3 = 8'b00000000;
 parameter INITREGBACKG_0_3 = 8'b00000000;
 
 parameter LOSE7 = 8'b10000001;
 parameter LOSE6 = 8'b01000100;
 parameter LOSE5 = 8'b00101000;
 parameter LOSE4 = 8'b00010000;
 parameter LOSE3 = 8'b00101000;
 parameter LOSE2 = 8'b01000100;
 parameter LOSE1 = 8'b10000010;
 parameter LOSE0 = 8'b11111111;
 
 parameter WIN7 = 8'b01111110;
 parameter WIN6 = 8'b10111101;
 parameter WIN5 = 8'b10111101;
 parameter WIN4 = 8'b01111110;
 parameter WIN3 = 8'b00011000;
 parameter WIN2 = 8'b00011000;
 parameter WIN1 = 8'b00111100;
 parameter WIN0 = 8'b01111110;
  
//=======================================================
//  PORT declarations
//=======================================================
output		[DISPLAY_DATAWIDTH-1:0] BB_SYSTEM_display_OutBUS;

output		BB_SYSTEM_max7219DIN_Out;
output		BB_SYSTEM_max7219NCS_Out;
output		BB_SYSTEM_max7219CLK_Out;

output 		BB_SYSTEM_startButton_Out;
output 		BB_SYSTEM_upButton_Out;
output 		BB_SYSTEM_downButton_Out;
output 		BB_SYSTEM_leftButton_Out;
output 		BB_SYSTEM_rightButton_Out;
output 		BB_SYSTEM_TEST0;
output 		BB_SYSTEM_TEST1;
output 		BB_SYSTEM_TEST2;

input		BB_SYSTEM_CLOCK_50;
input		BB_SYSTEM_RESET_InHigh;
input		BB_SYSTEM_startButton_InLow;
input		BB_SYSTEM_upButton_InLow;
input		BB_SYSTEM_downButton_InLow;
input		BB_SYSTEM_leftButton_InLow;
input		BB_SYSTEM_rightButton_InLow;
//=======================================================
//  REG/WIRE declarations
//=======================================================
wire  COLLISIONCOMPARATOR_EXIT_wire;
wire	[3:0]SC_STATEMACHINEPRINCIPAL_NEXTLEVEL_wire;
wire	[2:0]SC_STATEMACHINEPRINCIPAL_RESETLEVEL_wire;
wire	SC_STATEMACHINEPRINCIPAL_LIVEOUT_wire;
wire	SC_STATEMACHINEPRINCIPAL_LEVELOUT_wire;
wire	[7:0]SC_STATEMACHINEPRINCIPAL_LEVELOR_wire;
wire	[3:0]SC_LIVECOUNTER_data_OutBUS_wire;
wire	[3:0]SC_LEVELCOUNTER_data_OutBUS_wire;

// BUTTONs
wire 	BB_SYSTEM_startButton_InLow_cwire;
wire 	BB_SYSTEM_upButton_InLow_cwire;
wire 	BB_SYSTEM_downButton_InLow_cwire;
wire 	BB_SYSTEM_leftButton_InLow_cwire;
wire 	BB_SYSTEM_rightButton_InLow_cwire;

//POINT
wire	STATEMACHINEPOINT_clear_cwire;
wire	STATEMACHINEPOINT_load0_cwire;
wire	STATEMACHINEPOINT_load1_cwire;
wire	[1:0] STATEMACHINEPOINT_shiftselection_cwire;

wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data14_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data13_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data12_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data11_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data10_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data9_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data8_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data7_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data6_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data5_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data4_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data3_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data2_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data1_Out;
wire [DATAWIDTH_BUS-1:0] RegPOINTTYPE_2_POINTMATRIX_data0_Out;

//BACKGROUNG
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data14_Out;

wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data13_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data12_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data11_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data10_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data9_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data8_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data7_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data6_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data5_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data4_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data3_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data2_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data1_Out;
wire [DATAWIDTH_BUS-1:0] RegBACKGTYPE_2_BACKGMATRIX_data0_Out;

wire [7:0]DATA_FIXED_INITREGBACKG_0;
wire [7:0]DATA_FIXED_INITREGBACKG_1;
wire [7:0]DATA_FIXED_INITREGBACKG_2;
wire [7:0]DATA_FIXED_INITREGBACKG_3;
wire [7:0]DATA_FIXED_INITREGBACKG_4;
wire [7:0]DATA_FIXED_INITREGBACKG_5;
wire [7:0]DATA_FIXED_INITREGBACKG_6;
wire [7:0]DATA_FIXED_INITREGBACKG_7;
wire [7:0]DATA_FIXED_INITREGBACKG_8;
wire [7:0]DATA_FIXED_INITREGBACKG_9;
wire [7:0]DATA_FIXED_INITREGBACKG_10;
wire [7:0]DATA_FIXED_INITREGBACKG_11;
wire [7:0]DATA_FIXED_INITREGBACKG_12;wire [7:0]DATA_FIXED_INITREGBACKG_13;

wire [PRESCALER_DATAWIDTH-1:0] upSPEEDCOUNTER_data_BUS_wire;
wire SPEEDCOMPARATOR_2_STATEMACHINEBACKG_T0_cwire;
wire STATEMACHINEBACKG_clear_cwire;
wire STATEMACHINEBACKG_load_cwire;
wire [1:0] STATEMACHINEBACKG_shiftselection_cwire;
wire STATEMACHINEBACKG_upcount_cwire;

//BOTTOMSIDE COMPARATOR
wire BOTTOMSIDECOMPARATOR_2_STATEMACHINEBACKG_bottomside_cwire;

// GAME
wire [DATAWIDTH_BUS-1:0] regGAME_data7_wire;
wire [DATAWIDTH_BUS-1:0] regGAME_data6_wire;
wire [DATAWIDTH_BUS-1:0] regGAME_data5_wire;
wire [DATAWIDTH_BUS-1:0] regGAME_data4_wire;
wire [DATAWIDTH_BUS-1:0] regGAME_data3_wire;
wire [DATAWIDTH_BUS-1:0] regGAME_data2_wire;
wire [DATAWIDTH_BUS-1:0] regGAME_data1_wire;
wire [DATAWIDTH_BUS-1:0] regGAME_data0_wire;

wire 	[7:0] data_max;
wire 	[2:0] add;

wire [DATAWIDTH_BUS-1:0] upCOUNTER_2_BIN2BCD1_data_BUS_wire;
wire [DISPLAY_DATAWIDTH-1:0] BIN2BCD1_2_SEVENSEG1_data_BUS_wire;

//=======================================================
//  Structural coding
//=======================================================

//######################################################################
//#	INPUTS
//######################################################################
SC_DEBOUNCE1 SC_DEBOUNCE1_u0 (
// port map - connection between master ports and signals/registers   
	.SC_DEBOUNCE1_button_Out(BB_SYSTEM_startButton_InLow_cwire),
	.SC_DEBOUNCE1_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_DEBOUNCE1_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_DEBOUNCE1_button_In(~BB_SYSTEM_startButton_InLow)
);
SC_DEBOUNCE1 SC_DEBOUNCE1_u1 (
// port map - connection between master ports and signals/registers   
	.SC_DEBOUNCE1_button_Out(BB_SYSTEM_upButton_InLow_cwire),
	.SC_DEBOUNCE1_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_DEBOUNCE1_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_DEBOUNCE1_button_In(~BB_SYSTEM_upButton_InLow)
);
SC_DEBOUNCE1 SC_DEBOUNCE1_u2 (
// port map - connection between master ports and signals/registers   
	.SC_DEBOUNCE1_button_Out(BB_SYSTEM_downButton_InLow_cwire),
	.SC_DEBOUNCE1_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_DEBOUNCE1_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_DEBOUNCE1_button_In(~BB_SYSTEM_downButton_InLow)
);
SC_DEBOUNCE1 SC_DEBOUNCE1_u3 (
// port map - connection between master ports and signals/registers   
	.SC_DEBOUNCE1_button_Out(BB_SYSTEM_leftButton_InLow_cwire),
	.SC_DEBOUNCE1_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_DEBOUNCE1_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_DEBOUNCE1_button_In(~BB_SYSTEM_leftButton_InLow)
);
SC_DEBOUNCE1 SC_DEBOUNCE1_u4 (
// port map - connection between master ports and signals/registers   
	.SC_DEBOUNCE1_button_Out(BB_SYSTEM_rightButton_InLow_cwire),
	.SC_DEBOUNCE1_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_DEBOUNCE1_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_DEBOUNCE1_button_In(~BB_SYSTEM_rightButton_InLow)
);

//######################################################################
//#	POINT
//######################################################################
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_14)) SC_RegPOINTTYPE_u14 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data14_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data13_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data0_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_13)) SC_RegPOINTTYPE_u13 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data13_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data12_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data14_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_12)) SC_RegPOINTTYPE_u12 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data12_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data11_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data13_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_11)) SC_RegPOINTTYPE_u11 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data11_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data10_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data12_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_10)) SC_RegPOINTTYPE_u10 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data10_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data9_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data11_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_9)) SC_RegPOINTTYPE_u9 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data9_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data8_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data10_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_8)) SC_RegPOINTTYPE_u8 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data8_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data7_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data9_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_7)) SC_RegPOINTTYPE_u7 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data7_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data6_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data8_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_6)) SC_RegPOINTTYPE_u6 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data6_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data5_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data7_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_5)) SC_RegPOINTTYPE_u5 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data5_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data4_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data6_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_4)) SC_RegPOINTTYPE_u4 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data4_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data3_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data5_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_3)) SC_RegPOINTTYPE_u3 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data3_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data2_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data4_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_2)) SC_RegPOINTTYPE_u2 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data2_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data1_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data3_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_1)) SC_RegPOINTTYPE_u1 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data1_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data0_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data2_Out)
);
SC_RegPOINTTYPE #(.RegPOINTTYPE_DATAWIDTH(DATAWIDTH_BUS), .DATA_FIXED_INITREGPOINT(DATA_FIXED_INITREGPOINT_0)) SC_RegPOINTTYPE_u0 (
// port map - connection between master ports and signals/registers   
	.SC_RegPOINTTYPE_data_OutBUS(RegPOINTTYPE_2_POINTMATRIX_data0_Out),
	.SC_RegPOINTTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegPOINTTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegPOINTTYPE_clear_InLow(STATEMACHINEPOINT_clear_cwire),
	.SC_RegPOINTTYPE_load0_InLow(STATEMACHINEPOINT_load0_cwire),
	.SC_RegPOINTTYPE_load1_InLow(STATEMACHINEPOINT_load1_cwire),
	.SC_RegPOINTTYPE_shiftselection_In(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_RegPOINTTYPE_data0_InBUS(RegPOINTTYPE_2_POINTMATRIX_data14_Out),
	.SC_RegPOINTTYPE_data1_InBUS(RegPOINTTYPE_2_POINTMATRIX_data1_Out)
);

SC_STATEMACHINEPOINT SC_STATEMACHINEPOINT_u0 (
// port map - connection between master ports and signals/registers   
	.SC_STATEMACHINEPOINT_clear_OutLow(STATEMACHINEPOINT_clear_cwire), 
	.SC_STATEMACHINEPOINT_load0_OutLow(STATEMACHINEPOINT_load0_cwire), 
	.SC_STATEMACHINEPOINT_load1_OutLow(STATEMACHINEPOINT_load1_cwire), 
	.SC_STATEMACHINEPOINT_shiftselection_Out(STATEMACHINEPOINT_shiftselection_cwire),
	.SC_STATEMACHINEPOINT_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_STATEMACHINEPOINT_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_STATEMACHINEPOINT_startButton_InLow(BB_SYSTEM_startButton_InLow_cwire), 
	.SC_STATEMACHINEPOINT_upButton_InLow(BB_SYSTEM_upButton_InLow_cwire), 
	.SC_STATEMACHINEPOINT_downButton_InLow(BB_SYSTEM_downButton_InLow_cwire), 
	.SC_STATEMACHINEPOINT_leftButton_InLow(BB_SYSTEM_leftButton_InLow_cwire), 
	.SC_STATEMACHINEPOINT_rightButton_InLow(BB_SYSTEM_rightButton_InLow_cwire), 
	.SC_STATEMACHINEPOINT_bottomsidecomparator_InLow(BOTTOMSIDECOMPARATOR_2_STATEMACHINEBACKG_bottomside_cwire),
	.SC_STATEMACHINEPOINT_RESETLEVEL(SC_STATEMACHINEPRINCIPAL_RESETLEVEL_wire),
	.SC_STATEMACHINEPOINT_NEXTLEVEL(SC_STATEMACHINEPRINCIPAL_NEXTLEVEL_wire)
);

//######################################################################
//#	BACKGROUND
//######################################################################
SC_RegBACKTYPELAST SC_RegBACKTYPELAST_u14 (
// port map - connection between master ports and signals/registers   
	.SC_RegBACKTYPELAST_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data14_Out),
	.SC_RegBACKTYPELAST_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKTYPELAST_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKTYPELAST_NEXTLEVEL(SC_STATEMACHINEPRINCIPAL_NEXTLEVEL_wire),
	.SC_RegBACKTYPELAST_LEVELOR(SC_STATEMACHINEPRINCIPAL_LEVELOR_wire)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u13 (
// port map - connection between master ports and signals/registers 
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_13),  
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data13_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u12 (
// port map - connection between master ports and signals/registers 
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_12),  
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data12_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u11 (
// port map - connection between master ports and signals/registers 
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_11),  
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data11_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u10 (
// port map - connection between master ports and signals/registers
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_10),   
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data10_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u9 (
// port map - connection between master ports and signals/registers 
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_9),  
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data9_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u8 (
// port map - connection between master ports and signals/registers
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_8),   
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data8_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u7 (
// port map - connection between master ports and signals/registers
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_7),   
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data7_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u6 (
// port map - connection between master ports and signals/registers
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_6),   
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data6_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u5 (
// port map - connection between master ports and signals/registers 
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_5),  
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data5_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u4 (
// port map - connection between master ports and signals/registers 
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_4),  
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data4_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u3 (
// port map - connection between master ports and signals/registers
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_3),   
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data3_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u2 (
// port map - connection between master ports and signals/registers 
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_2),  
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data2_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u1 (
// port map - connection between master ports and signals/registers
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_1),   
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data1_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_RegBACKGTYPE #(.RegBACKGTYPE_DATAWIDTH(DATAWIDTH_BUS)) SC_RegBACKGTYPE_u0 (
// port map - connection between master ports and signals/registers
	.DATA_FIXED_INITREGBACKG(DATA_FIXED_INITREGBACKG_0),
	.SC_RegBACKGTYPE_data_OutBUS(RegBACKGTYPE_2_BACKGMATRIX_data0_Out),
	.SC_RegBACKGTYPE_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_RegBACKGTYPE_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_RegBACKGTYPE_clear_InLow(STATEMACHINEBACKG_clear_cwire),	
	.SC_RegBACKGTYPE_load_InLow(STATEMACHINEBACKG_load_cwire),
	.SC_RegBACKGTYPE_shiftselection_In(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_RegBACKGTYPE_data_InBUS(DATA_FIXED_INITREGBACKG_0)
);
SC_STATEMACHINEBACKG SC_STATEMACHINEBACKG_u0 (
// port map - connection between master ports and signals/registers   
	.SC_STATEMACHINEBACKG_clear_OutLow(STATEMACHINEBACKG_clear_cwire), 
	.SC_STATEMACHINEBACKG_load_OutLow(STATEMACHINEBACKG_load_cwire), 
	.SC_STATEMACHINEBACKG_shiftselection_Out(STATEMACHINEBACKG_shiftselection_cwire),
	.SC_STATEMACHINEBACKG_upcount_out(STATEMACHINEBACKG_upcount_cwire),
	.SC_STATEMACHINEBACKG_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_STATEMACHINEBACKG_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_STATEMACHINEBACKG_startButton_InLow(BB_SYSTEM_startButton_InLow_cwire),
	.SC_STATEMACHINEBACKG_T0_InLow(SPEEDCOMPARATOR_2_STATEMACHINEBACKG_T0_cwire)
);

SC_STATEMACHINEPRINCIPAL SC_STATEMACHINEPRINCIPAL_u0 (   
	.SC_STATEMACHINEPRINCIPAL_NEXTLEVEL(SC_STATEMACHINEPRINCIPAL_NEXTLEVEL_wire), 
	.SC_STATEMACHINEPRINCIPAL_RESETLEVEL(SC_STATEMACHINEPRINCIPAL_RESETLEVEL_wire), 
	.SC_STATEMACHINEPRINCIPAL_LIVEOUT(SC_STATEMACHINEPRINCIPAL_LIVEOUT_wire),
	.SC_STATEMACHINEPRINCIPAL_LEVELOUT(SC_STATEMACHINEPRINCIPAL_LEVELOUT_wire),
	.SC_STATEMACHINEPRINCIPAL_LEVELOR(SC_STATEMACHINEPRINCIPAL_LEVELOR_wire),
	.SC_STATEMACHINEPRINCIPAL_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_STATEMACHINEPRINCIPAL_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_STATEMACHINEPRINCIPAL_HOUSES(RegBACKGTYPE_2_BACKGMATRIX_data14_Out),
	.SC_STATEMACHINEPRINCIPAL_CEXIT(COLLISIONCOMPARATOR_EXIT_wire),
	.SC_STATEMACHINEPRINCIPAL_LIVECOUNT(SC_LIVECOUNTER_data_OutBUS_wire),
	.SC_STATEMACHINEPRINCIPAL_LEVELCOUNT(SC_LEVELCOUNTER_data_OutBUS_wire)
);
//#SPEED
SC_upSPEEDCOUNTER #(.upSPEEDCOUNTER_DATAWIDTH(PRESCALER_DATAWIDTH)) SC_upSPEEDCOUNTER_u0 (
// port map - connection between master ports and signals/registers   
	.SC_upSPEEDCOUNTER_data_OutBUS(upSPEEDCOUNTER_data_BUS_wire),
	.SC_upSPEEDCOUNTER_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_upSPEEDCOUNTER_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_upSPEEDCOUNTER_upcount_InLow(STATEMACHINEBACKG_upcount_cwire)
);

CC_SPEEDCOMPARATOR #(.SPEEDCOMPARATOR_DATAWIDTH(PRESCALER_DATAWIDTH)) CC_SPEEDCOMPARATOR_u0 (
	.CC_SPEEDCOMPARATOR_T0_OutLow(SPEEDCOMPARATOR_2_STATEMACHINEBACKG_T0_cwire),
	.CC_SPEEDCOMPARATOR_data_InBUS(upSPEEDCOUNTER_data_BUS_wire)
);

SC_LIVECOUNTER SC_LIVECOUNTER_u0 (  
	.SC_LIVECOUNTER_data_OutBUS(SC_LIVECOUNTER_data_OutBUS_wire),
	.SC_LIVECOUNTER_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_LIVECOUNTER_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_LIVECOUNTER_CUENTA(SC_STATEMACHINEPRINCIPAL_LIVEOUT_wire)
);

SC_LEVELCOUNTER SC_LEVELCOUNTER_u0 (  
	.SC_LEVELCOUNTER_data_OutBUS(SC_LEVELCOUNTER_data_OutBUS_wire),
	.SC_LEVELCOUNTER_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_LEVELCOUNTER_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_LEVELCOUNTER_CUENTA(SC_STATEMACHINEPRINCIPAL_LEVELOUT_wire)
);
//######################################################################
//#	COMPARATOR END OF MATRIX (BOTTON SIDE)
//######################################################################
CC_BOTTOMSIDECOMPARATOR #(.BOTTOMSIDECOMPARATOR_DATAWIDTH(DATAWIDTH_BUS)) CC_BOTTOMSIDECOMPARATOR_u0 (
	.CC_BOTTOMSIDECOMPARATOR_bottomside_OutLow(BOTTOMSIDECOMPARATOR_2_STATEMACHINEBACKG_bottomside_cwire),
	.CC_BOTTOMSIDECOMPARATOR_data_InBUS(RegPOINTTYPE_2_POINTMATRIX_data0_Out)
);

//######################################################################
//#	COMPARATOR SCREEN
//######################################################################
CC_SCREENCOMPARATOR CC_SCREENCOMPARATOR_u0 (
	.CC_SCREENCOMPARATOR_0(regGAME_data0_wire),
	.CC_SCREENCOMPARATOR_1(regGAME_data1_wire),
	.CC_SCREENCOMPARATOR_2(regGAME_data2_wire),
	.CC_SCREENCOMPARATOR_3(regGAME_data3_wire),
	.CC_SCREENCOMPARATOR_4(regGAME_data4_wire),
	.CC_SCREENCOMPARATOR_5(regGAME_data5_wire),
	.CC_SCREENCOMPARATOR_6(regGAME_data6_wire),
	.CC_SCREENCOMPARATOR_7(regGAME_data7_wire),

	.CC_SCREENCOMPARATOR_POINT_0(RegPOINTTYPE_2_POINTMATRIX_data0_Out),
	.CC_SCREENCOMPARATOR_POINT_1(RegPOINTTYPE_2_POINTMATRIX_data1_Out),
	.CC_SCREENCOMPARATOR_POINT_2(RegPOINTTYPE_2_POINTMATRIX_data2_Out),
	.CC_SCREENCOMPARATOR_POINT_3(RegPOINTTYPE_2_POINTMATRIX_data3_Out),
	.CC_SCREENCOMPARATOR_POINT_4(RegPOINTTYPE_2_POINTMATRIX_data4_Out),
	.CC_SCREENCOMPARATOR_POINT_5(RegPOINTTYPE_2_POINTMATRIX_data5_Out),
	.CC_SCREENCOMPARATOR_POINT_6(RegPOINTTYPE_2_POINTMATRIX_data6_Out),
	.CC_SCREENCOMPARATOR_POINT_7(RegPOINTTYPE_2_POINTMATRIX_data7_Out),
	.CC_SCREENCOMPARATOR_POINT_8(RegPOINTTYPE_2_POINTMATRIX_data8_Out),
	.CC_SCREENCOMPARATOR_POINT_9(RegPOINTTYPE_2_POINTMATRIX_data9_Out),
	.CC_SCREENCOMPARATOR_POINT_10(RegPOINTTYPE_2_POINTMATRIX_data10_Out),
	.CC_SCREENCOMPARATOR_POINT_11(RegPOINTTYPE_2_POINTMATRIX_data11_Out),
	.CC_SCREENCOMPARATOR_POINT_12(RegPOINTTYPE_2_POINTMATRIX_data12_Out),
	.CC_SCREENCOMPARATOR_POINT_13(RegPOINTTYPE_2_POINTMATRIX_data13_Out),
	.CC_SCREENCOMPARATOR_POINT_14(RegPOINTTYPE_2_POINTMATRIX_data14_Out),
	
	.CC_SCREENCOMPARATOR_BACK_0(RegBACKGTYPE_2_BACKGMATRIX_data0_Out),
	.CC_SCREENCOMPARATOR_BACK_1(RegBACKGTYPE_2_BACKGMATRIX_data1_Out),
	.CC_SCREENCOMPARATOR_BACK_2(RegBACKGTYPE_2_BACKGMATRIX_data2_Out),
	.CC_SCREENCOMPARATOR_BACK_3(RegBACKGTYPE_2_BACKGMATRIX_data3_Out),
	.CC_SCREENCOMPARATOR_BACK_4(RegBACKGTYPE_2_BACKGMATRIX_data4_Out),
	.CC_SCREENCOMPARATOR_BACK_5(RegBACKGTYPE_2_BACKGMATRIX_data5_Out),
	.CC_SCREENCOMPARATOR_BACK_6(RegBACKGTYPE_2_BACKGMATRIX_data6_Out),
	.CC_SCREENCOMPARATOR_BACK_7(RegBACKGTYPE_2_BACKGMATRIX_data7_Out),
	.CC_SCREENCOMPARATOR_BACK_8(RegBACKGTYPE_2_BACKGMATRIX_data8_Out),
	.CC_SCREENCOMPARATOR_BACK_9(RegBACKGTYPE_2_BACKGMATRIX_data9_Out),
	.CC_SCREENCOMPARATOR_BACK_10(RegBACKGTYPE_2_BACKGMATRIX_data10_Out),
	.CC_SCREENCOMPARATOR_BACK_11(RegBACKGTYPE_2_BACKGMATRIX_data11_Out),
	.CC_SCREENCOMPARATOR_BACK_12(RegBACKGTYPE_2_BACKGMATRIX_data12_Out),
	.CC_SCREENCOMPARATOR_BACK_13(RegBACKGTYPE_2_BACKGMATRIX_data13_Out),
	.CC_SCREENCOMPARATOR_BACK_14(RegBACKGTYPE_2_BACKGMATRIX_data14_Out),
	
	.CC_SCREENCOMPARATOR_LOSE_0(LOSE0),
	.CC_SCREENCOMPARATOR_LOSE_1(LOSE1),
	.CC_SCREENCOMPARATOR_LOSE_2(LOSE2),
	.CC_SCREENCOMPARATOR_LOSE_3(LOSE3),
	.CC_SCREENCOMPARATOR_LOSE_4(LOSE4),
	.CC_SCREENCOMPARATOR_LOSE_5(LOSE5),
	.CC_SCREENCOMPARATOR_LOSE_6(LOSE6),
	.CC_SCREENCOMPARATOR_LOSE_7(LOSE7),
	
	.CC_SCREENCOMPARATOR_WIN_0(WIN0),
	.CC_SCREENCOMPARATOR_WIN_1(WIN1),
	.CC_SCREENCOMPARATOR_WIN_2(WIN2),
	.CC_SCREENCOMPARATOR_WIN_3(WIN3),
	.CC_SCREENCOMPARATOR_WIN_4(WIN4),
	.CC_SCREENCOMPARATOR_WIN_5(WIN5),
	.CC_SCREENCOMPARATOR_WIN_6(WIN6),
	.CC_SCREENCOMPARATOR_WIN_7(WIN7),
	
	.CC_SCREENCOMPARATOR_LOSE(SC_STATEMACHINEPRINCIPAL_RESETLEVEL_wire),
	.CC_SCREENCOMPARATOR_WIN(SC_STATEMACHINEPRINCIPAL_NEXTLEVEL_wire)
);
//######################################################################
//#	COMPARATOR COLLISION
//######################################################################
CC_COLLISIONCOMPARATOR CC_COLLISIONCOMPARATOR_u0 (
	.CC_COLLISIONCOMPARATOR_EXIT(COLLISIONCOMPARATOR_EXIT_wire),

	.CC_COLLISIONCOMPARATOR_POINT_0(RegPOINTTYPE_2_POINTMATRIX_data0_Out),
	.CC_COLLISIONCOMPARATOR_POINT_1(RegPOINTTYPE_2_POINTMATRIX_data1_Out),
	.CC_COLLISIONCOMPARATOR_POINT_2(RegPOINTTYPE_2_POINTMATRIX_data2_Out),
	.CC_COLLISIONCOMPARATOR_POINT_3(RegPOINTTYPE_2_POINTMATRIX_data3_Out),
	.CC_COLLISIONCOMPARATOR_POINT_4(RegPOINTTYPE_2_POINTMATRIX_data4_Out),
	.CC_COLLISIONCOMPARATOR_POINT_5(RegPOINTTYPE_2_POINTMATRIX_data5_Out),
	.CC_COLLISIONCOMPARATOR_POINT_6(RegPOINTTYPE_2_POINTMATRIX_data6_Out),
	.CC_COLLISIONCOMPARATOR_POINT_7(RegPOINTTYPE_2_POINTMATRIX_data7_Out),
	.CC_COLLISIONCOMPARATOR_POINT_8(RegPOINTTYPE_2_POINTMATRIX_data8_Out),
	.CC_COLLISIONCOMPARATOR_POINT_9(RegPOINTTYPE_2_POINTMATRIX_data9_Out),
	.CC_COLLISIONCOMPARATOR_POINT_10(RegPOINTTYPE_2_POINTMATRIX_data10_Out),
	.CC_COLLISIONCOMPARATOR_POINT_11(RegPOINTTYPE_2_POINTMATRIX_data11_Out),
	.CC_COLLISIONCOMPARATOR_POINT_12(RegPOINTTYPE_2_POINTMATRIX_data12_Out),
	.CC_COLLISIONCOMPARATOR_POINT_13(RegPOINTTYPE_2_POINTMATRIX_data13_Out),
	.CC_COLLISIONCOMPARATOR_POINT_14(RegPOINTTYPE_2_POINTMATRIX_data14_Out),
	
	.CC_COLLISIONCOMPARATOR_BACK_0(RegBACKGTYPE_2_BACKGMATRIX_data0_Out),
	.CC_COLLISIONCOMPARATOR_BACK_1(RegBACKGTYPE_2_BACKGMATRIX_data1_Out),
	.CC_COLLISIONCOMPARATOR_BACK_2(RegBACKGTYPE_2_BACKGMATRIX_data2_Out),
	.CC_COLLISIONCOMPARATOR_BACK_3(RegBACKGTYPE_2_BACKGMATRIX_data3_Out),
	.CC_COLLISIONCOMPARATOR_BACK_4(RegBACKGTYPE_2_BACKGMATRIX_data4_Out),
	.CC_COLLISIONCOMPARATOR_BACK_5(RegBACKGTYPE_2_BACKGMATRIX_data5_Out),
	.CC_COLLISIONCOMPARATOR_BACK_6(RegBACKGTYPE_2_BACKGMATRIX_data6_Out),
	.CC_COLLISIONCOMPARATOR_BACK_7(RegBACKGTYPE_2_BACKGMATRIX_data7_Out),
	.CC_COLLISIONCOMPARATOR_BACK_8(RegBACKGTYPE_2_BACKGMATRIX_data8_Out),
	.CC_COLLISIONCOMPARATOR_BACK_9(RegBACKGTYPE_2_BACKGMATRIX_data9_Out),
	.CC_COLLISIONCOMPARATOR_BACK_10(RegBACKGTYPE_2_BACKGMATRIX_data10_Out),
	.CC_COLLISIONCOMPARATOR_BACK_11(RegBACKGTYPE_2_BACKGMATRIX_data11_Out),
	.CC_COLLISIONCOMPARATOR_BACK_12(RegBACKGTYPE_2_BACKGMATRIX_data12_Out),
	.CC_COLLISIONCOMPARATOR_BACK_13(RegBACKGTYPE_2_BACKGMATRIX_data13_Out),
	.CC_COLLISIONCOMPARATOR_BACK_14(RegBACKGTYPE_2_BACKGMATRIX_data14_Out),
	
	.CC_COLLISIONCOMPARATOR_LOSE(SC_STATEMACHINEPRINCIPAL_RESETLEVEL_wire),
	.CC_COLLISIONCOMPARATOR_WIN(SC_STATEMACHINEPRINCIPAL_NEXTLEVEL_wire)
);
//######################################################################
//#	COMPARATOR LEVEL
//######################################################################
CC_LEVELCOMPARATOR CC_LEVELCOMPARATOR_u0(
	.CC_SCREEN_0(DATA_FIXED_INITREGBACKG_0),
	.CC_SCREEN_1(DATA_FIXED_INITREGBACKG_1),
	.CC_SCREEN_2(DATA_FIXED_INITREGBACKG_2),
	.CC_SCREEN_3(DATA_FIXED_INITREGBACKG_3),
	.CC_SCREEN_4(DATA_FIXED_INITREGBACKG_4),
	.CC_SCREEN_5(DATA_FIXED_INITREGBACKG_5),
	.CC_SCREEN_6(DATA_FIXED_INITREGBACKG_6),
	.CC_SCREEN_7(DATA_FIXED_INITREGBACKG_7),
	.CC_SCREEN_8(DATA_FIXED_INITREGBACKG_8),
	.CC_SCREEN_9(DATA_FIXED_INITREGBACKG_9),
	.CC_SCREEN_10(DATA_FIXED_INITREGBACKG_10),
	.CC_SCREEN_11(DATA_FIXED_INITREGBACKG_11),
	.CC_SCREEN_12(DATA_FIXED_INITREGBACKG_12),
	.CC_SCREEN_13(DATA_FIXED_INITREGBACKG_13),

	.CC_LEVELCOMPARATOR_LEVELCOUNTER(SC_LEVELCOUNTER_data_OutBUS_wire)
);
//######################################################################
//#	TO LED MATRIZ: VISUALIZATION
//######################################################################
assign data_max =(add==3'b000)?{regGAME_data0_wire[7],regGAME_data1_wire[7],regGAME_data2_wire[7],regGAME_data3_wire[7],regGAME_data4_wire[7],regGAME_data5_wire[7],regGAME_data6_wire[7],regGAME_data7_wire[7]}:
	       (add==3'b001)?{regGAME_data0_wire[6],regGAME_data1_wire[6],regGAME_data2_wire[6],regGAME_data3_wire[6],regGAME_data4_wire[6],regGAME_data5_wire[6],regGAME_data6_wire[6],regGAME_data7_wire[6]}:
	       (add==3'b010)?{regGAME_data0_wire[5],regGAME_data1_wire[5],regGAME_data2_wire[5],regGAME_data3_wire[5],regGAME_data4_wire[5],regGAME_data5_wire[5],regGAME_data6_wire[5],regGAME_data7_wire[5]}:
	       (add==3'b011)?{regGAME_data0_wire[4],regGAME_data1_wire[4],regGAME_data2_wire[4],regGAME_data3_wire[4],regGAME_data4_wire[4],regGAME_data5_wire[4],regGAME_data6_wire[4],regGAME_data7_wire[4]}:
	       (add==3'b100)?{regGAME_data0_wire[3],regGAME_data1_wire[3],regGAME_data2_wire[3],regGAME_data3_wire[3],regGAME_data4_wire[3],regGAME_data5_wire[3],regGAME_data6_wire[3],regGAME_data7_wire[3]}:
	       (add==3'b101)?{regGAME_data0_wire[2],regGAME_data1_wire[2],regGAME_data2_wire[2],regGAME_data3_wire[2],regGAME_data4_wire[2],regGAME_data5_wire[2],regGAME_data6_wire[2],regGAME_data7_wire[2]}:
	       (add==3'b110)?{regGAME_data0_wire[1],regGAME_data1_wire[1],regGAME_data2_wire[1],regGAME_data3_wire[1],regGAME_data4_wire[1],regGAME_data5_wire[1],regGAME_data6_wire[1],regGAME_data7_wire[1]}:
						{regGAME_data0_wire[0],regGAME_data1_wire[0],regGAME_data2_wire[0],regGAME_data3_wire[0],regGAME_data4_wire[0],regGAME_data5_wire[0],regGAME_data6_wire[0],regGAME_data7_wire[0]};
									 
matrix_ctrl matrix_ctrl_unit_0( 
.max7219_din(BB_SYSTEM_max7219DIN_Out),//max7219_din 
.max7219_ncs(BB_SYSTEM_max7219NCS_Out),//max7219_ncs 
.max7219_clk(BB_SYSTEM_max7219CLK_Out),//max7219_clk
.disp_data(data_max), 
.disp_addr(add),
.intensity(4'hA),
.clk(BB_SYSTEM_CLOCK_50),
.reset(BB_SYSTEM_RESET_InHigh) //~lowRst_System
 ); 
 
//~ imagen img1(
//~ .act_add(add), 
//~ .max_in(data_max) );

//~ SC_CTRLMATRIX SC_CTRLMATRIX_u0( 
//~ .SC_CTRLMATRIX_max7219DIN_Out(BB_SYSTEM_max7219DIN_Out),	//max7219_din 
//~ .SC_CTRLMATRIX_max7219NCS_out(BB_SYSTEM_max7219NCS_Out),	//max7219_ncs 
//~ .SC_CTRLMATRIX_max7219CLK_Out(BB_SYSTEM_max7219CLK_Out),	//max7219_clk
//~ .SC_CTRLMATRIX_dispdata(data_max), 
//~ .SC_CTRLMATRIX_dispaddr(add),
//~ .SC_CTRLMATRIX_intensity(4'hA),
//~ .SC_CTRLMATRIX_CLOCK_50(BB_SYSTEM_CLOCK_50),
//~ .SC_CTRLMATRIX_RESET_InHigh(~BB_SYSTEM_RESET_InHigh) 		//~lowRst_System
 //~ ); 
 
//~ SC_IMAGE SC_IMAGE_u0(
//~ .SC_IMAGE_actadd(add), 
//~ .SC_IMAGE_maxin(data_max) );

//######################################################################
//#	TO TEST
//######################################################################

assign BB_SYSTEM_startButton_Out = BB_SYSTEM_startButton_InLow_cwire;
assign BB_SYSTEM_upButton_Out = BB_SYSTEM_upButton_InLow_cwire;
assign BB_SYSTEM_downButton_Out = BB_SYSTEM_downButton_InLow_cwire;
assign BB_SYSTEM_leftButton_Out = BB_SYSTEM_leftButton_InLow_cwire;
assign BB_SYSTEM_rightButton_Out = BB_SYSTEM_rightButton_InLow_cwire;
//TO TEST
assign BB_SYSTEM_TEST0 = BB_SYSTEM_startButton_InLow_cwire;
assign BB_SYSTEM_TEST1 = BB_SYSTEM_startButton_InLow_cwire;
assign BB_SYSTEM_TEST2 = BB_SYSTEM_startButton_InLow_cwire;

//######################################################################
//#	TO 7SEG
//######################################################################

CC_BIN2BCD1 CC_BIN2BCD1_u0 (
// port map - connection between master ports and signals/registers   
	.CC_BIN2BCD_bcd_OutBUS(BIN2BCD1_2_SEVENSEG1_data_BUS_wire),
	.CC_BIN2BCD_bin_InBUS(upCOUNTER_2_BIN2BCD1_data_BUS_wire)
);

CC_SEVENSEG1 CC_SEVENSEG1_u0 (
// port map - connection between master ports and signals/registers   
	.CC_SEVENSEG1_an(BB_SYSTEM_display_OutBUS[11:8]),
	.CC_SEVENSEG1_a(BB_SYSTEM_display_OutBUS[0]),
	.CC_SEVENSEG1_b(BB_SYSTEM_display_OutBUS[1]),
	.CC_SEVENSEG1_c(BB_SYSTEM_display_OutBUS[2]),
	.CC_SEVENSEG1_d(BB_SYSTEM_display_OutBUS[3]),
	.CC_SEVENSEG1_e(BB_SYSTEM_display_OutBUS[4]),
	.CC_SEVENSEG1_f(BB_SYSTEM_display_OutBUS[5]),
	.CC_SEVENSEG1_g(BB_SYSTEM_display_OutBUS[6]),
	.CC_SEVENSEG1_dp(BB_SYSTEM_display_OutBUS[7]),
	.CC_SEVENSEG1_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.CC_SEVENSEG1_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.CC_SEVENSEG1_in0(BIN2BCD1_2_SEVENSEG1_data_BUS_wire[3:0]),
	.CC_SEVENSEG1_in1(BIN2BCD1_2_SEVENSEG1_data_BUS_wire[7:4]),
	.CC_SEVENSEG1_in2(BIN2BCD1_2_SEVENSEG1_data_BUS_wire[11:8]),
	.CC_SEVENSEG1_in3(BIN2BCD1_2_SEVENSEG1_data_BUS_wire[11:8])
);

SC_upCOUNTER #(.upCOUNTER_DATAWIDTH(DATAWIDTH_BUS)) SC_upCOUNTER_u0 (
// port map - connection between master ports and signals/registers   
	.SC_upCOUNTER_data_OutBUS(upCOUNTER_2_BIN2BCD1_data_BUS_wire),
	.SC_upCOUNTER_CLOCK_50(BB_SYSTEM_CLOCK_50),
	.SC_upCOUNTER_RESET_InHigh(BB_SYSTEM_RESET_InHigh),
	.SC_upCOUNTER_upcount_InLow(STATEMACHINEPOINT_load0_cwire)
);

endmodule
